module top_module ( input a, input b, output out );
    mod_a g1(a,b,out);
    	

endmodule
